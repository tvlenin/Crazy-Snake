`timescale 1ns / 1ps

module Random_Generator(
	input clock,
	input [5:0] yValues,
	input [5:0] xValues
);

endmodule
