`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:54:20 04/25/2017 
// Design Name: 
// Module Name:    font_rom 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module font_rom(
    input clk,
    input [10:0] addr,
    output [7:0] data
    );
	 reg [10:0] addr_reg;
	 always@(posedge clk)
		addr_reg <= addr;
	
	 always@*
		case(addr_reg)
			//espacio vacio
			11'h000: data = 8'b00000000;
			11'h03a: data = 8'b00000000;
			11'h002: data = 8'b00000000;
			11'h003: data = 8'b00000000;
			11'h004: data = 8'b00000000;
			11'h005: data = 8'b00000000;
			11'h006: data = 8'b00000000;
			11'h007: data = 8'b00000000;
			11'h008: data = 8'b00000000;
			11'h009: data = 8'b00000000;
			11'h00a: data = 8'b00000000;
			11'h00b: data = 8'b00000000;
			11'h00c: data = 8'b00000000;
			11'h00d: data = 8'b00000000;
			11'h00f: data = 8'b00000000;

			11'h010: data =8'b00000000;//  0
			11'h011: data =8'b00000000;//  1
			11'h012: data =8'b00010000;//  2    *
			11'h013: data =8'b00111000;//  3   ***
			11'h014: data =8'b01101100;//  4  ** **
			11'h015: data =8'b11000110;//  5 **   **
			11'h016: data =8'b11000110;//  6 **   **
			11'h017: data =8'b11111110;//  7 *******
			11'h018: data =8'b11000110;//  8 **   **
			11'h019: data =8'b11000110;//  9 **   **
			11'h01a: data =8'b11000110;//  a **   **
			11'h01b: data =8'b11000110;//  b **   **
			11'h01c: data =8'b00000000;//  c
			11'h01d: data =8'b00000000;//  d
			11'h01e: data =8'b00000000;//  e
			11'h01f: data =8'b00000000;//  f


			11'h020: data =8'b00000000;//   1
			11'h021: data =8'b11111100;//   2 ******
			11'h022: data =8'b01100110;//   3  **  **
			11'h023: data =8'b01100110;//   4  **  **
			11'h024: data =8'b01100110;//   5  **  **
			11'h025: data =8'b01111100;//   6  *****
			11'h026: data =8'b01100110;//   7  **  **
			11'h027: data =8'b01100110;//   8  **  **
			11'h028: data =8'b01100110;//   9  **  **
			11'h029: data =8'b01100110;//   a  **  **
			11'h02a: data =8'b11111100;//   b ******
			11'h02b: data =8'b00000000;//   c
			11'h02c: data =8'b00000000;//   d
			11'h02d: data =8'b00000000;//   e
			11'h02f: data =8'b00000000;//   f
			//C: code x43
			11'h030: data =8'b00000000;//   0
			11'h031: data =8'b00000000;//   1
			11'h032: data =8'b00111100;//   2   ****
			11'h033: data =8'b01100110;//   3  **  **
			11'h034: data =8'b11000010;//   4 **    *
			11'h035: data =8'b11000000;//   5 **
			11'h036: data =8'b11000000;//   6 **
			11'h037: data =8'b11000000;//   7 **
			11'h038: data =8'b11000000;//   8 **
			11'h039: data =8'b11000010;//   9 **    *
			11'h03a: data =8'b01100110;//   a  **  **
			11'h03b: data =8'b00111100;//   b   ****
			11'h03c: data =8'b00000000;//   c
			11'h03d: data =8'b00000000;//   d
			11'h03e: data =8'b00000000;//   e
			11'h03f: data =8'b00000000;//   f
			//D: code x44
			11'h040: data =8'b00000000;//   0
			11'h041: data =8'b00000000;//   1
			11'h042: data =8'b11111000;//   2 *****
			11'h043: data =8'b01101100;//   3  ** **
			11'h044: data =8'b01100110;//   4  **  **
			11'h045: data =8'b01100110;//   5  **  **
			11'h046: data =8'b01100110;//   6  **  **
			11'h047: data =8'b01100110;//   7  **  **
			11'h048: data =8'b01100110;//   8  **  **
			11'h049: data =8'b01100110;//   9  **  **
			11'h04a: data =8'b01101100;//   a  ** **
			11'h04b: data =8'b11111000;//   b *****
			11'h04c: data =8'b00000000;//   c
			11'h04d: data =8'b00000000;//   d
			11'h04e: data =8'b00000000;//   e
			11'h04f: data =8'b00000000;//   f
			//code x45
			11'h050: data =8'b00000000;//   0
			11'h051: data =8'b00000000;//   1
			11'h052: data =8'b11111110;//   2 *******
			11'h053: data =8'b01100110;//   3  **  **
			11'h054: data =8'b01100010;//   4  **   *
			11'h055: data =8'b01101000;//   5  ** *
			11'h056: data =8'b01111000;//   6  ****
			11'h057: data =8'b01101000;//   7  ** *
			11'h058: data =8'b01100000;//   8  **
			11'h059: data =8'b01100010;//   9  **   *
			11'h05a: data =8'b01100110;//   a  **  **
			11'h05b: data =8'b11111110;//   b *******
			11'h05c: data =8'b00000000;//   c
			11'h05d: data =8'b00000000;//   d
			11'h05e: data =8'b00000000;//   e
			11'h05f: data =8'b00000000;//   f
			//code x46
			11'h060: data =8'b00000000;//   0
			11'h061: data =8'b00000000;//   1
			11'h062: data =8'b11111110;//   2 *******
			11'h063: data =8'b01100110;//   3  **  **
			11'h064: data =8'b01100010;//   4  **   *
			11'h065: data =8'b01101000;//   5  ** *
			11'h066: data =8'b01111000;//   6  ****
			11'h067: data =8'b01101000;//   7  ** *
			11'h068: data =8'b01100000;//   8  **
			11'h069: data =8'b01100000;//   9  **
			11'h06a: data =8'b01100000;//   a  **
			11'h06b: data =8'b11110000;//   b ****
			11'h06c: data =8'b00000000;//   c
			11'h06d: data =8'b00000000;//   d
			11'h06e: data =8'b00000000;//   e
			11'h06f: data =8'b00000000;//   f
			//code x47
			11'h070: data =8'b00000000;//   0
			11'h071: data =8'b00000000;//   1
			11'h072: data =8'b00111100;//   2   ****
			11'h073: data =8'b01100110;//   3  **  **
			11'h074: data =8'b11000010;//   4 **    *
			11'h075: data =8'b11000000;//   5 **
			11'h076: data =8'b11000000;//   6 **
			11'h077: data =8'b11011110;//   7 ** ****
			11'h078: data =8'b11000110;//   8 **   **
			11'h079: data =8'b11000110;//   9 **   **
			11'h07a: data =8'b01100110;//   a  **  **
			11'h07b: data =8'b00111010;//   b   *** *
			11'h07c: data =8'b00000000;//   c
			11'h07d: data =8'b00000000;//   d
			11'h07e: data =8'b00000000;//   e
			11'h07f: data =8'b00000000;//   f
			//H: code x48
			11'h080: data =8'b00000000;//   0
			11'h081: data =8'b00000000;//   1
			11'h082: data =8'b11000110;//   2 **   **
			11'h083: data =8'b11000110;//   3 **   **
			11'h084: data =8'b11000110;//   4 **   **
			11'h085: data =8'b11000110;//   5 **   **
			11'h086: data =8'b11111110;//   6 *******
			11'h087: data =8'b11000110;//   7 **   **
			11'h088: data =8'b11000110;//   8 **   **
			11'h089: data =8'b11000110;//   9 **   **
			11'h08a: data =8'b11000110;//   a **   **
			11'h08b: data =8'b11000110;//   b **   **
			11'h08c: data =8'b00000000;//   c
			11'h08d: data =8'b00000000;//   d
			11'h08e: data =8'b00000000;//   e
			11'h08f: data =8'b00000000;//   f
			//I: code x49
			11'h090: data =8'b00000000;//   0
			11'h091: data =8'b00000000;//   1
			11'h091: data =8'b00111100;//   2   ****
			11'h091: data =8'b00011000;//   3    **
			11'h091: data =8'b00011000;//   4    **
			11'h091: data =8'b00011000;//   5    **
			11'h091: data =8'b00011000;//   6    **
			11'h091: data =8'b00011000;//   7    **
			11'h091: data =8'b00011000;//   8    **
			11'h091: data =8'b00011000;//   9    **
			11'h091: data =8'b00011000;//   a    **
			11'h091: data =8'b00111100;//   b   ****
			11'h091: data =8'b00000000;//   c
			11'h091: data =8'b00000000;//   d
			11'h091: data =8'b00000000;//   e
			11'h091: data =8'b00000000;//   f
			//J: code x4a
			11'h100: data =8'b00000000;//   0
			11'h101: data =8'b00000000;//   1
			11'h102: data =8'b00011110;//   2    ****
			11'h103: data =8'b00001100;//   3     **
			11'h104: data =8'b00001100;//   4     **
			11'h105: data =8'b00001100;//   5     **
			11'h106: data =8'b00001100;//   6     **
			11'h107: data =8'b00001100;//   7     **
			11'h108: data =8'b11001100;//   8 **  **
			11'h109: data =8'b11001100;//   9 **  **
			11'h10a: data =8'b11001100;//   a **  **
			11'h10b: data =8'b01111000;//   b  ****
			11'h10c: data =8'b00000000;//   c
			11'h10d: data =8'b00000000;//   d
			11'h10e: data =8'b00000000;//   e
			11'h10f: data =8'b00000000;//   f
			//K: code x4b
			11'h110: data =8'b00000000;//   0
			11'h111: data =8'b00000000;//   1
			11'h112: data =8'b11100110;//   2 ***  **
			11'h113: data =8'b01100110;//   3  **  **
			11'h114: data =8'b01100110;//   4  **  **
			11'h115: data =8'b01101100;//   5  ** **
			11'h116: data =8'b01111000;//   6  ****
			11'h117: data =8'b01111000;//   7  ****
			11'h118: data =8'b01101100;//   8  ** **
			11'h119: data =8'b01100110;//   9  **  **
			11'h11a: data =8'b01100110;//   a  **  **
			11'h11b: data =8'b11100110;//   b ***  **
			11'h11c: data =8'b00000000;//   c
			11'h11d: data =8'b00000000;//   d
			11'h11e: data =8'b00000000;//   e
			11'h11f: data =8'b00000000;//   f
			//L: code x4c
			11'h120: data =8'b00000000;//   0
			11'h121: data =8'b00000000;//   1
			11'h122: data =8'b11110000;//   2 ****
			11'h123: data =8'b01100000;//   3  **
			11'h124: data =8'b01100000;//   4  **
			11'h125: data =8'b01100000;//   5  **
			11'h126: data =8'b01100000;//   6  **
			11'h127: data =8'b01100000;//   7  **
			11'h128: data =8'b01100000;//   8  **
			11'h129: data =8'b01100010;//   9  **   *
			11'h12a: data =8'b01100110;//   a  **  **
			11'h12b: data =8'b11111110;//   b *******
			11'h12c: data =8'b00000000;//   c
			11'h12d: data =8'b00000000;//   d
			11'h12e: data =8'b00000000;//   e
			11'h12f: data =8'b00000000;//   f
			//M: code x4d
			11'h130: data =8'b00000000;//   0
			11'h131: data =8'b00000000;//   1
			11'h132: data =8'b11000011;//   2 **    **
			11'h133: data =8'b11100111;//   3 ***  ***
			11'h134: data =8'b11111111;//   4 ********
			11'h135: data =8'b11111111;//   5 ********
			11'h136: data =8'b11011011;//   6 ** ** **
			11'h137: data =8'b11000011;//   7 **    **
			11'h138: data =8'b11000011;//   8 **    **
			11'h139: data =8'b11000011;//   9 **    **
			11'h13a: data =8'b11000011;//   a **    **
			11'h13b: data =8'b11000011;//   b **    **
			11'h13c: data =8'b00000000;//   c
			11'h13d: data =8'b00000000;//   d
			11'h13e: data =8'b00000000;//   e
			11'h13f: data =8'b00000000;//   f
			//N: code x4e
			11'h140: data =8'b00000000;//   0
			11'h141: data =8'b00000000;//   1
			11'h142: data =8'b11000110;//   2 **   **
			11'h143: data =8'b11100110;//   3 ***  **
			11'h144: data =8'b11110110;//   4 **** **
			11'h145: data =8'b11111110;//   5 *******
			11'h146: data =8'b11011110;//   6 ** ****
			11'h147: data =8'b11001110;//   7 **  ***
			11'h148: data =8'b11000110;//   8 **   **
			11'h149: data =8'b11000110;//   9 **   **
			11'h14a: data =8'b11000110;//   a **   **
			11'h14b: data =8'b11000110;//   b **   **
			11'h14c: data =8'b00000000;//   c
			11'h14d: data =8'b00000000;//   d
			11'h14e: data =8'b00000000;//   e
			11'h14f: data =8'b00000000;//   f
			//O: code x4f
			11'h150: data =8'b00000000;//   0
			11'h151: data =8'b00000000;//   1
			11'h152: data =8'b01111100;//   2  *****
			11'h153: data =8'b11000110;//   3 **   **
			11'h154: data =8'b11000110;//   4 **   **
			11'h155: data =8'b11000110;//   5 **   **
			11'h156: data =8'b11000110;//   6 **   **
			11'h157: data =8'b11000110;//   7 **   **
			11'h158: data =8'b11000110;//   8 **   **
			11'h159: data =8'b11000110;//   9 **   **
			11'h15a: data =8'b11000110;//   a **   **
			11'h15b: data =8'b01111100;//   b  *****
			11'h15c: data =8'b00000000;//   c
			11'h15d: data =8'b00000000;//   d
			11'h15e: data =8'b00000000;//   e
			11'h15f: data =8'b00000000;//   f
			//P: code x50
			11'h160: data =8'b00000000;//   0
			11'h161: data =8'b00000000;//   1
			11'h162: data =8'b11111100;//   2 ******
			11'h163: data =8'b01100110;//   3  **  **
			11'h164: data =8'b01100110;//   4  **  **
			11'h165: data =8'b01100110;//   5  **  **
			11'h166: data =8'b01111100;//   6  *****
			11'h167: data =8'b01100000;//   7  **
			11'h168: data =8'b01100000;//   8  **
			11'h169: data =8'b01100000;//   9  **
			11'h16a: data =8'b01100000;//   a  **
			11'h16b: data =8'b11110000;//   b ****
			11'h16c: data =8'b00000000;//   c
			11'h16d: data =8'b00000000;//   d
			11'h16e: data =8'b00000000;//   e
			11'h16f: data =8'b00000000;//   f
			//Q: code x510
			11'h170: data =8'b00000000;//   0
			11'h171: data =8'b00000000;//   1
			11'h172: data =8'b01111100;//   2  *****
			11'h173: data =8'b11000110;//   3 **   **
			11'h174: data =8'b11000110;//   4 **   **
			11'h175: data =8'b11000110;//   5 **   **
			11'h176: data =8'b11000110;//   6 **   **
			11'h177: data =8'b11000110;//   7 **   **
			11'h178: data =8'b11000110;//   8 **   **
			11'h179: data =8'b11010110;//   9 ** * **
			11'h17a: data =8'b11011110;//   a ** ****
			11'h17b: data =8'b01111100;//   b  *****
			11'h17c: data =8'b00001100;//   c     **
			11'h17d: data =8'b00001110;//   d     ***
			11'h17e: data =8'b00000000;//   e
			11'h17f: data =8'b00000000;//   f
			//code x52
			11'h180: data =8'b00000000;//   0
			11'h181: data =8'b00000000;//   1
			11'h182: data =8'b11111100;//   2 ******
			11'h183: data =8'b01100110;//   3  **  **
			11'h184: data =8'b01100110;//   4  **  **
			11'h185: data =8'b01100110;//   5  **  **
			11'h186: data =8'b01111100;//   6  *****
			11'h187: data =8'b01101100;//   7  ** **
			11'h188: data =8'b01100110;//   8  **  **
			11'h189: data =8'b01100110;//   9  **  **
			11'h18a: data =8'b01100110;//   a  **  **
			11'h18b: data =8'b11100110;//   b ***  **
			11'h18c: data =8'b00000000;//   c
			11'h18d: data =8'b00000000;//   d
			11'h18e: data =8'b00000000;//   e
			11'h18f: data =8'b00000000;//   f
			//code x53
			11'h190: data =8'b00000000;//   0
			11'h191: data =8'b00000000;//   1
			11'h192: data =8'b01111100;//   2  *****
			11'h193: data =8'b11000110;//   3 **   **
			11'h194: data =8'b11000110;//   4 **   **
			11'h195: data =8'b01100000;//   5  **
			11'h196: data =8'b00111000;//   6   ***
			11'h197: data =8'b00001100;//   7     **
			11'h198: data =8'b00000110;//   8      **
			11'h199: data =8'b11000110;//   9 **   **
			11'h19a: data =8'b11000110;//   a **   **
			11'h19b: data =8'b01111100;//   b  *****
			11'h19c: data =8'b00000000;//   c
			11'h19d: data =8'b00000000;//   d
			11'h19e: data =8'b00000000;//   e
			11'h19f: data =8'b00000000;//   f
			//code x54
			11'h200: data =8'b00000000;//   0
			11'h201: data =8'b00000000;//   1
			11'h202: data =8'b11111111;//   2 ********
			11'h203: data =8'b11011011;//   3 ** ** **
			11'h204: data =8'b10011001;//   4 *  **  *
			11'h205: data =8'b00011000;//   5    **
			11'h206: data =8'b00011000;//   6    **
			11'h207: data =8'b00011000;//   7    **
			11'h208: data =8'b00011000;//   8    **
			11'h209: data =8'b00011000;//   9    **
			11'h20a: data =8'b00011000;//   a    **
			11'h20b: data =8'b00111100;//   b   ****
			11'h20c: data =8'b00000000;//   c
			11'h20d: data =8'b00000000;//   d
			11'h20e: data =8'b00000000;//   e
			11'h20f: data =8'b00000000;//   f
			//code x55
			11'h210: data =8'b00000000;//   0
			11'h211: data =8'b00000000;//   1
			11'h212: data =8'b11000110;//   2 **   **
			11'h213: data =8'b11000110;//   3 **   **
			11'h214: data =8'b11000110;//   4 **   **
			11'h215: data =8'b11000110;//   5 **   **
			11'h216: data =8'b11000110;//   6 **   **
			11'h217: data =8'b11000110;//   7 **   **
			11'h218: data =8'b11000110;//   8 **   **
			11'h219: data =8'b11000110;//   9 **   **
			11'h21a: data =8'b11000110;//   a **   **
			11'h21b: data =8'b01111100;//   b  *****
			11'h21c: data =8'b00000000;//   c
			11'h21d: data =8'b00000000;//   d
			11'h21e: data =8'b00000000;//   e
			11'h21f: data =8'b00000000;//   f
			//code x56
			11'h220: data =8'b00000000;//   0
			11'h221: data =8'b00000000;//   1
			11'h222: data =8'b11000011;//   2 **    **
			11'h223: data =8'b11000011;//   3 **    **
			11'h224: data =8'b11000011;//   4 **    **
			11'h225: data =8'b11000011;//   5 **    **
			11'h226: data =8'b11000011;//   6 **    **
			11'h227: data =8'b11000011;//   7 **    **
			11'h228: data =8'b11000011;//   8 **    **
			11'h229: data =8'b01100110;//   9  **  **
			11'h22a: data =8'b00111100;//   a   ****
			11'h22b: data =8'b00011000;//   b    **
			11'h22c: data =8'b00000000;//   c
			11'h22d: data =8'b00000000;//   d
			11'h22e: data =8'b00000000;//   e
			11'h22f: data =8'b00000000;//   f
			//code x57
			11'h230: data =8'b00000000;//   0
			11'h231: data =8'b00000000;//   1
			11'h232: data =8'b11000011;//   2 **    **
			11'h233: data =8'b11000011;//   3 **    **
			11'h234: data =8'b11000011;//   4 **    **
			11'h235: data =8'b11000011;//   5 **    **
			11'h236: data =8'b11000011;//   6 **    **
			11'h237: data =8'b11011011;//   7 ** ** **
			11'h238: data =8'b11011011;//   8 ** ** **
			11'h239: data =8'b11111111;//   9 ********
			11'h23a: data =8'b01100110;//   a  **  **
			11'h23b: data =8'b01100110;//   b  **  **
			11'h23c: data =8'b00000000;//   c
			11'h23d: data =8'b00000000;//   d
			11'h23e: data =8'b00000000;//   e
			11'h23f: data =8'b00000000;//   f

			//code x58
			11'h240: data =8'b00000000;//   0
			11'h241: data =8'b00000000;//   1
			11'h242: data =8'b11000011;//   2 **    **
			11'h243: data =8'b11000011;//   3 **    **
			11'h244: data =8'b01100110;//   4  **  **
			11'h245: data =8'b00111100;//   5   ****
			11'h246: data =8'b00011000;//   6    **
			11'h247: data =8'b00011000;//   7    **
			11'h248: data =8'b00111100;//   8   ****
			11'h249: data =8'b01100110;//   9  **  **
			11'h24a: data =8'b11000011;//   a **    **
			11'h24b: data =8'b11000011;//   b **    **
			11'h24c: data =8'b00000000;//   c
			11'h24d: data =8'b00000000;//   d
			11'h24e: data =8'b00000000;//   e
			11'h24f: data =8'b00000000;//   f
			//code x59
			11'h250: data =8'b00000000;//   0
			11'h251: data =8'b00000000;//   1
			11'h252: data =8'b11000011;//   2 **    **
			11'h253: data =8'b11000011;//   3 **    **
			11'h254: data =8'b11000011;//   4 **    **
			11'h255: data =8'b01100110;//   5  **  **
			11'h256: data =8'b00111100;//   6   ****
			11'h257: data =8'b00011000;//   7    **
			11'h258: data =8'b00011000;//   8    **
			11'h259: data =8'b00011000;//   9    **
			11'h25a: data =8'b00011000;//   a    **
			11'h25b: data =8'b00111100;//   b   ****
			11'h25c: data =8'b00000000;//   c
			11'h25d: data =8'b00000000;//   d
			11'h25e: data =8'b00000000;//   e
			11'h25f: data =8'b00000000;//   f
			//code x5a
			11'h260: data =8'b00000000;//   0
			11'h261: data =8'b00000000;//   1
			11'h262: data =8'b11111111;//   2 ********
			11'h263: data =8'b11000011;//   3 **    **
			11'h264: data =8'b10000110;//   4 *    **
			11'h265: data =8'b00001100;//   5     **
			11'h266: data =8'b00011000;//   6    **
			11'h267: data =8'b00110000;//   7   **
			11'h268: data =8'b01100000;//   8  **
			11'h269: data =8'b11000001;//   9 **     *
			11'h26a: data =8'b11000011;//   a **    **
			11'h26b: data =8'b11111111;//   b ********
			11'h26c: data =8'b00000000;//   c
			11'h26d: data =8'b00000000;//   d
			11'h26e: data =8'b00000000;//   e
			11'h26f: data =8'b00000000;//   f

	 
		endcase

endmodule
